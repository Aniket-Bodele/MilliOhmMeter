CircuitMaker Text
5.6
Probes: 1
U1_6
Transient Analysis
0 585 178 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
220 60 30 120 10
176 80 1534 803
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
56 C:\Users\Dell\OneDrive\Desktop\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 1702 537
9961490 0
0
6 Title:
5 Name:
0
0
0
27
13 Var Resistor~
219 801 268 0 3 7
0 23 4 3
0
0 0 848 90
8 100k 25%
8 -4 64 4
3 R11
25 -14 46 -6
0
0
32 %DA %1 %2 25000
%DB %2 %3 75000
0
0
4 SIP3
7

0 1 2 3 1 2 3 0
82 0 0 512 1 0 0 0
1 R
5130 0 0
2
5.90072e-315 0
0
11 Multimeter~
205 619 93 0 21 21
0 6 24 25 5 0 0 0 0 0
32 53 48 48 46 48 109 65 0 0
0 86
0
0 0 16464 270
6 1.000u
-21 -19 21 -11
3 MM2
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
391 0 0
2
5.90072e-315 0
0
11 Multimeter~
205 567 321 0 21 21
0 9 26 27 8 0 0 0 0 0
32 53 48 48 46 48 109 65 0 0
0 86
0
0 0 16464 270
6 1.000u
-21 -19 21 -11
3 MM1
-11 -29 10 -21
0
0
28 R1%D %1 %2 %V
%D %2 %4 DC 0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.90072e-315 0
0
11 Multimeter~
205 1013 255 0 21 21
0 7 28 29 2 0 0 0 0 0
32 52 46 56 57 57 32 86 0 0
0 82
0
0 0 16464 0
8 100.0Meg
-28 -19 28 -11
3 MM0
-11 -29 10 -21
0
0
11 %D %1 %4 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
1 R
3421 0 0
2
5.90072e-315 0
0
2 +V
167 698 154 0 1 3
0 16
0
0 0 54256 512
3 10V
-11 -22 10 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.90072e-315 0
0
2 +V
167 699 209 0 1 3
0 15
0
0 0 54256 180
4 -10V
3 -2 31 6
2 V8
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5572 0 0
2
5.90072e-315 0
0
2 +V
167 702 347 0 1 3
0 17
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8901 0 0
2
5.90072e-315 0
0
2 +V
167 708 408 0 1 3
0 14
0
0 0 54256 180
4 -10V
3 -2 31 6
2 V6
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.90072e-315 0
0
2 +V
167 900 262 0 1 3
0 11
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4747 0 0
2
5.90072e-315 0
0
2 +V
167 902 325 0 1 3
0 10
0
0 0 54256 180
3 10V
6 -2 27 6
2 V4
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
972 0 0
2
5.90072e-315 0
0
2 +V
167 531 185 0 1 3
0 13
0
0 0 54256 0
2 9V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3472 0 0
2
5.90072e-315 0
0
2 +V
167 533 252 0 1 3
0 12
0
0 0 54256 180
3 -9V
6 -2 27 6
2 V2
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9998 0 0
2
5.90072e-315 0
0
7 Ground~
168 995 172 0 1 3
0 2
0
0 0 53360 90
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3536 0 0
2
5.90072e-315 0
0
7 Ground~
168 587 290 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4597 0 0
2
5.90072e-315 0
0
8 Op-Amp5~
219 901 292 0 5 11
0 20 18 11 10 7
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U4
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3835 0 0
2
5.90072e-315 0
0
8 Op-Amp5~
219 703 371 0 5 11
0 22 4 17 14 19
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U3
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
3670 0 0
2
5.90072e-315 0
0
2 +V
167 502 384 0 1 3
0 8
0
0 0 54256 180
3 -9V
6 -2 27 6
2 V1
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
5.90072e-315 0
0
8 Op-Amp5~
219 697 177 0 5 11
0 6 3 16 15 21
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U2
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
9323 0 0
2
5.90072e-315 0
0
8 Op-Amp5~
219 530 215 0 5 11
0 22 2 13 12 6
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U1
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
317 0 0
2
5.90072e-315 0
0
9 Resistor~
219 833 374 0 2 5
0 18 19
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
5.90072e-315 0
0
9 Resistor~
219 944 318 0 2 5
0 18 7
0
0 0 880 90
2 1k
8 0 22 8
2 R8
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4299 0 0
2
5.90072e-315 0
0
9 Resistor~
219 904 173 0 3 5
0 2 20 -1
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
5.90072e-315 0
0
9 Resistor~
219 807 176 0 2 5
0 20 21
0
0 0 880 180
2 1k
-7 -14 7 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7876 0 0
2
5.90072e-315 0
0
9 Resistor~
219 742 341 0 2 5
0 19 4
0
0 0 880 90
4 330k
2 0 30 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6369 0 0
2
5.90072e-315 0
0
9 Resistor~
219 753 197 0 2 5
0 3 21
0
0 0 880 90
4 330k
2 0 30 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9172 0 0
2
5.90072e-315 0
0
9 Resistor~
219 505 304 0 2 5
0 9 22
0
0 0 880 90
2 18
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7100 0 0
2
5.90072e-315 0
0
9 Resistor~
219 594 251 0 2 5
0 22 5
0
0 0 880 90
1 1
12 0 19 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3820 0 0
2
5.90072e-315 0
0
37
0 1 3 0 0 4096 0 0 25 28 0 3
752 225
752 215
753 215
2 0 4 0 0 12416 0 1 0 0 0 4
793 266
793 288
804 288
804 312
0 0 4 0 0 8192 0 0 0 2 29 9
804 308
809 308
809 348
804 348
804 350
776 350
776 315
748 315
748 321
1 0 3 0 0 0 0 25 0 0 28 3
753 215
753 220
752 220
4 2 5 0 0 4224 0 2 27 0 0 3
603 125
603 233
594 233
0 1 6 0 0 4224 0 0 2 33 0 3
585 215
585 75
603 75
0 1 7 0 0 4224 0 0 4 24 0 3
944 292
988 292
988 278
0 4 2 0 0 8192 0 0 4 26 0 6
973 173
973 210
1066 210
1066 288
1038 288
1038 278
4 1 8 0 0 4224 0 3 17 0 0 3
551 353
502 353
502 369
1 1 9 0 0 8320 0 26 3 0 0 5
505 322
505 326
543 326
543 303
551 303
4 1 10 0 0 8320 0 15 10 0 0 3
901 305
902 305
902 310
3 1 11 0 0 8320 0 15 9 0 0 3
901 279
900 279
900 271
1 4 12 0 0 4224 0 12 19 0 0 3
533 237
533 228
530 228
1 3 13 0 0 8320 0 11 19 0 0 3
531 194
530 194
530 202
1 4 14 0 0 4224 0 8 16 0 0 3
708 393
708 384
703 384
1 4 15 0 0 8320 0 6 18 0 0 3
699 194
697 194
697 190
1 4 15 0 0 0 0 6 18 0 0 3
699 194
697 194
697 190
3 1 16 0 0 4224 0 18 5 0 0 3
697 164
697 163
698 163
1 3 17 0 0 4224 0 7 16 0 0 3
702 356
702 358
703 358
1 3 16 0 0 0 0 5 18 0 0 3
698 163
698 164
697 164
1 0 18 0 0 4096 0 20 0 0 23 2
851 374
883 374
0 2 19 0 0 8320 0 0 20 30 0 3
753 371
753 374
815 374
2 1 18 0 0 4224 0 15 21 0 0 4
883 286
883 374
944 374
944 336
5 2 7 0 0 0 0 15 21 0 0 3
919 292
944 292
944 300
0 1 20 0 0 4224 0 0 15 27 0 3
851 176
851 298
883 298
1 1 2 0 0 0 0 22 13 0 0 2
922 173
988 173
1 2 20 0 0 0 0 23 22 0 0 3
825 176
886 176
886 173
2 3 3 0 0 12416 0 18 1 0 0 7
679 171
655 171
655 225
761 225
761 208
805 208
805 246
2 2 4 0 0 8320 0 16 24 0 0 6
685 365
685 321
748 321
748 321
742 321
742 323
1 5 19 0 0 0 0 24 16 0 0 5
742 359
742 371
753 371
753 371
721 371
0 2 21 0 0 8192 0 0 25 32 0 3
751 176
753 176
753 179
5 2 21 0 0 8320 0 18 23 0 0 3
715 177
715 176
789 176
5 1 6 0 0 0 0 19 18 0 0 3
548 215
679 215
679 183
1 1 22 0 0 8320 0 27 16 0 0 4
594 269
647 269
647 377
685 377
1 2 2 0 0 4224 0 14 19 0 0 4
587 284
458 284
458 209
512 209
0 2 22 0 0 0 0 0 26 37 0 3
512 269
505 269
505 286
1 1 22 0 0 0 0 27 19 0 0 3
594 269
512 269
512 221
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
